module orTest(result, a ,b);
input[4:0] a,b;
output[4:0] result;


assign result = a | b;

endmodule