library verilog;
use verilog.vl_types.all;
entity mips_testbench is
end mips_testbench;
